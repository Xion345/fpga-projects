../../library/basic/counter_mod_m.vhd