../../library/uart/uart_rxtx_clock.vhd