../../library/vga/vga_tiles.vhd