../../library/uart/uart_rx.vhd