../../library/uart/uart_dma.vhd