../../library/block_ram/block_ram.vhd