../../library/uart/uart_tx.vhd