../../library/vga/vga_sync.vhd